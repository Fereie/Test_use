module counter_8b
input a
input b

and o,a,b

